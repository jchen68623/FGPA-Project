`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Team Members: Carlos Perez, Ramos Jiuru Chen
//
// Control Signals:
//		EX: ALUSrc, ALUOp, RegDst
//		M: Branch, MemRead, MemWrite, Zero
//		PCSrc
//		WB: RegWrite, MemtoReg
//		 ALUSrcTop(shift select)
//
////////////////////////////////////////////////////////////////////////////////

module ID_EX_reg(
// inputs
Reset,
Hi, Lo,
Clock, PCadder, ALUSrc, RegDst, RegWrite, MemRead, MemWrite, MemtoReg, Branch, ALUop, ReadData1, ReadData2,
instruction15_0, instruction20_16, instruction15_11, mthi, mtlo, WriteEnable, ReadEnable, DataWidth, jumpAddress, jumpSrc,jregSrc, LinkStoreSel,
Rs, Rt, ControlWrite,
// outputs
PCadder_out, ALUSrc_out, RegDst_out, RegWrite_out, MemRead_out, MemWrite_out, MemtoReg_out, Branch_out, ALUop_out, ReadData1_out, ReadData2_out, 
instruction15_0_out, instruction20_16_out, instruction15_11_out, mthi_out, mtlo_out, WriteEnable_out, ReadEnable_out, DataWidth_out, jumpAddress_out, jumpSrc_out, jregSrc_out, LinkStoreSel_out,
Hi_out, Lo_out,
Rs_out, Rt_out
);
	//::INPUTS::
	input Clock;
	input Reset;
	input [31:0] PCadder;
	
	// Control signals generated by controller
	input ALUSrc, RegWrite, MemRead, MemWrite, MemtoReg, Branch;
	input [1:0] RegDst;
	input [5:0] ALUop;
	input [1:0] DataWidth;
	
	// two register values read from the register file
	input [31:0] ReadData1;
	input [31:0] ReadData2;
	
	// potential destination registers (Rd I[15:0] and I[20-16])
	input [31:0] instruction15_0;
	input [4:0] instruction20_16;
	input [4:0] instruction15_11;
	
	input mthi, mtlo, WriteEnable, ReadEnable;
	
	input [31:0] jumpAddress;
	input jumpSrc;
	input jregSrc;
	input LinkStoreSel;
	input [4:0] Rs, Rt;
	output reg [4:0] Rs_out, Rt_out;
	
	input ControlWrite;
	//::OUTPUTS::
	output reg [31:0]  PCadder_out;
	
	// Control signals
	output reg ALUSrc_out, RegWrite_out, MemRead_out, MemWrite_out, MemtoReg_out, Branch_out;
	output reg [1:0] RegDst_out;
	output reg [5:0] ALUop_out;
	output reg [1:0] DataWidth_out;
	
	// two register values read from the register file
	output reg [31:0] ReadData1_out;
	output reg [31:0] ReadData2_out;
	
	// sign extended offset field
//	output reg [31:0] signExtend_out; // offset[31:16] + instruction[15:0] renamed to instruction15_0_out
	
	// potential destination registers (Rd I[15:0] and I[20-16])
	output reg [31:0] instruction15_0_out;
	output reg [4:0] instruction20_16_out, instruction15_11_out;
	
	output reg mthi_out, mtlo_out, WriteEnable_out, ReadEnable_out;
	
	output reg [31:0] jumpAddress_out;
	output reg jumpSrc_out;
	output reg jregSrc_out;
	output reg LinkStoreSel_out;
	
	input [31:0] Hi;
	input [31:0] Lo;
	output reg [31:0] Hi_out;
	output reg [31:0] Lo_out;
	
	// zero outputs initially
	initial begin
		PCadder_out <= 0;
		ALUSrc_out <= 0;
		RegDst_out <= 0;
		RegWrite_out <= 0;
		MemRead_out <= 0;
		MemWrite_out <= 0;
		MemtoReg_out <= 0;
		Branch_out <= 0;
		//ALUSrcTop_out <= 0;
		ALUop_out <= 0;
		DataWidth_out <= 0;
		ReadData1_out <= 0;
		ReadData2_out <= 0;
		instruction15_0_out <= 0;
		instruction20_16_out <= 0;
		instruction15_11_out <= 0;
		mthi_out <= 0;
		mtlo_out <= 0;
		WriteEnable_out <= 0;
		ReadEnable_out <= 0;
		jumpAddress_out <= 0;
		Hi_out <= 0;
		Lo_out <= 0;
		jumpSrc_out <= 0;
		jregSrc_out <= 0;
		LinkStoreSel_out <= 0;
		Rs_out <= 0;
		Rt_out <= 0;
	end
	
//	always @(*) begin
//	   if (Reset == 1) begin
//            PCadder_out <= 0;
//            ALUSrc_out <= 0;
//            RegDst_out <= 0;
//            RegWrite_out <= 0;
//            MemRead_out <= 0;
//            MemWrite_out <= 0;
//            MemtoReg_out <= 0;
//            Branch_out <= 0;
//            //ALUSrcTop_out <= 0;
//            ALUop_out <= 0;
//            DataWidth_out <= 0;
//            ReadData1_out <= 0;
//            ReadData2_out <= 0;
//            instruction15_0_out <= 0;
//            instruction20_16_out <= 0;
//            instruction15_11_out <= 0;
//            mthi_out <= 0;
//            mtlo_out <= 0;
//            WriteEnable_out <= 0;
//            ReadEnable_out <= 0;
//            jumpAddress_out <= 0;
//            Hi_out <= 0;
//            Lo_out <= 0;
//            jumpSrc_out <= 0;
//            jregSrc_out <= 0;
//            LinkStoreSel_out <= 0;
//            Rs_out <= 0;
//            Rt_out <= 0;	   
//	   end
//	end
	
	always @(posedge Clock) begin
	    if (Reset == 1) begin
             PCadder_out <= 0;
             ALUSrc_out <= 0;
             RegDst_out <= 0;
             RegWrite_out <= 0;
             MemRead_out <= 0;
             MemWrite_out <= 0;
             MemtoReg_out <= 0;
             Branch_out <= 0;
             //ALUSrcTop_out <= 0;
             ALUop_out <= 0;
             DataWidth_out <= 0;
             ReadData1_out <= 0;
             ReadData2_out <= 0;
             instruction15_0_out <= 0;
             instruction20_16_out <= 0;
             instruction15_11_out <= 0;
             mthi_out <= 0;
             mtlo_out <= 0;
             WriteEnable_out <= 0;
             ReadEnable_out <= 0;
             jumpAddress_out <= 0;
             Hi_out <= 0;
             Lo_out <= 0;
             jumpSrc_out <= 0;
             jregSrc_out <= 0;
             LinkStoreSel_out <= 0;
             Rs_out <= 0;
             Rt_out <= 0;       
        end
        
        if (ControlWrite == 0) begin
            PCadder_out <= 0;
            ALUSrc_out <= 0;
            RegDst_out <= 0;
            RegWrite_out <= 0;
            MemRead_out <= 0;
            MemWrite_out <= 0;
            MemtoReg_out <= 0;
            Branch_out <= 0;
            //ALUSrcTop_out <= 0;
            ALUop_out <= 0;
            DataWidth_out <= 0;
            ReadData1_out <= 0;
            ReadData2_out <= 0;
            instruction15_0_out <= 0;
            instruction20_16_out <= 0;
            instruction15_11_out <= 0;
            mthi_out <= 0;
            mtlo_out <= 0;
            WriteEnable_out <= 0;
            ReadEnable_out <= 0;
            jumpAddress_out <= 0;
            Hi_out <= 0;
            Lo_out <= 0;
            jumpSrc_out <= 0;
            jregSrc_out <= 0;
            LinkStoreSel_out <= 0;
            Rs_out <= 0;
            Rt_out <= 0;
        end
        
        else if (ControlWrite == 1) begin
            PCadder_out <= PCadder;
            ALUSrc_out <= ALUSrc;
            RegDst_out <= RegDst;
            RegWrite_out <= RegWrite;
            MemRead_out <= MemRead;
            MemWrite_out <= MemWrite;
            MemtoReg_out <= MemtoReg;
            Branch_out <= Branch;
            //ALUSrcTop_out <= ALUSrcTop;
            ALUop_out <= ALUop;
            DataWidth_out <= DataWidth;
            ReadData1_out <= ReadData1;
            ReadData2_out <= ReadData2;
            instruction15_0_out <= instruction15_0;
            instruction20_16_out <= instruction20_16;
            instruction15_11_out <= instruction15_11;
            mthi_out <= mthi;
            mtlo_out <= mtlo;
            WriteEnable_out <= WriteEnable;
            ReadEnable_out <= ReadEnable;
            jumpAddress_out <= jumpAddress;
            jumpSrc_out <= jumpSrc;
            jregSrc_out <= jregSrc;
            LinkStoreSel_out <= LinkStoreSel;
            Hi_out <= Hi;
            Lo_out <= Lo;
            Rs_out <= Rs;
            Rt_out <= Rt;
        end
    end
    
endmodule